module leastALU();








endmodule
