module mux_2x1_32bit(a, b, s, r);

	input [31:0]a;
	input [31:0]b; 
	input s;
	output [31:0]r;
	
	
	// r = s'a + sb
	
	
	



endmodule
